module h;    
initial begin $display("Hello World"); $finish; end

	endmodule
